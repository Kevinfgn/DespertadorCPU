// DespertadorCPU_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DespertadorCPU_tb (
	);

	wire        despertadorcpu_inst_clk_bfm_clk_clk;              // DespertadorCPU_inst_clk_bfm:clk -> [DespertadorCPU_inst:clk_clk, DespertadorCPU_inst_reset_bfm:clk]
	wire  [0:0] despertadorcpu_inst_btnapagar_bfm_conduit_export; // DespertadorCPU_inst_btnapagar_bfm:sig_export -> DespertadorCPU_inst:btnapagar_export
	wire  [0:0] despertadorcpu_inst_btnhora_bfm_conduit_export;   // DespertadorCPU_inst_btnhora_bfm:sig_export -> DespertadorCPU_inst:btnhora_export
	wire  [0:0] despertadorcpu_inst_btnmin_bfm_conduit_export;    // DespertadorCPU_inst_btnmin_bfm:sig_export -> DespertadorCPU_inst:btnmin_export
	wire        despertadorcpu_inst_buzzer_export;                // DespertadorCPU_inst:buzzer_export -> DespertadorCPU_inst_buzzer_bfm:sig_export
	wire  [6:0] despertadorcpu_inst_hora1_export;                 // DespertadorCPU_inst:hora1_export -> DespertadorCPU_inst_hora1_bfm:sig_export
	wire  [6:0] despertadorcpu_inst_hora2_export;                 // DespertadorCPU_inst:hora2_export -> DespertadorCPU_inst_hora2_bfm:sig_export
	wire  [6:0] despertadorcpu_inst_min1_export;                  // DespertadorCPU_inst:min1_export -> DespertadorCPU_inst_min1_bfm:sig_export
	wire  [6:0] despertadorcpu_inst_min2_export;                  // DespertadorCPU_inst:min2_export -> DespertadorCPU_inst_min2_bfm:sig_export
	wire  [0:0] despertadorcpu_inst_swinicio_bfm_conduit_export;  // DespertadorCPU_inst_swinicio_bfm:sig_export -> DespertadorCPU_inst:swinicio_export
	wire  [0:0] despertadorcpu_inst_swmodo_bfm_conduit_export;    // DespertadorCPU_inst_swmodo_bfm:sig_export -> DespertadorCPU_inst:swmodo_export
	wire        despertadorcpu_inst_reset_bfm_reset_reset;        // DespertadorCPU_inst_reset_bfm:reset -> DespertadorCPU_inst:reset_reset_n

	DespertadorCPU despertadorcpu_inst (
		.btnapagar_export (despertadorcpu_inst_btnapagar_bfm_conduit_export), // btnapagar.export
		.btnhora_export   (despertadorcpu_inst_btnhora_bfm_conduit_export),   //   btnhora.export
		.btnmin_export    (despertadorcpu_inst_btnmin_bfm_conduit_export),    //    btnmin.export
		.buzzer_export    (despertadorcpu_inst_buzzer_export),                //    buzzer.export
		.clk_clk          (despertadorcpu_inst_clk_bfm_clk_clk),              //       clk.clk
		.hora1_export     (despertadorcpu_inst_hora1_export),                 //     hora1.export
		.hora2_export     (despertadorcpu_inst_hora2_export),                 //     hora2.export
		.min1_export      (despertadorcpu_inst_min1_export),                  //      min1.export
		.min2_export      (despertadorcpu_inst_min2_export),                  //      min2.export
		.reset_reset_n    (despertadorcpu_inst_reset_bfm_reset_reset),        //     reset.reset_n
		.swinicio_export  (despertadorcpu_inst_swinicio_bfm_conduit_export),  //  swinicio.export
		.swmodo_export    (despertadorcpu_inst_swmodo_bfm_conduit_export)     //    swmodo.export
	);

	altera_conduit_bfm despertadorcpu_inst_btnapagar_bfm (
		.sig_export (despertadorcpu_inst_btnapagar_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm despertadorcpu_inst_btnhora_bfm (
		.sig_export (despertadorcpu_inst_btnhora_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm despertadorcpu_inst_btnmin_bfm (
		.sig_export (despertadorcpu_inst_btnmin_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 despertadorcpu_inst_buzzer_bfm (
		.sig_export (despertadorcpu_inst_buzzer_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) despertadorcpu_inst_clk_bfm (
		.clk (despertadorcpu_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0003 despertadorcpu_inst_hora1_bfm (
		.sig_export (despertadorcpu_inst_hora1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 despertadorcpu_inst_hora2_bfm (
		.sig_export (despertadorcpu_inst_hora2_export)  // conduit.export
	);

	altera_conduit_bfm_0003 despertadorcpu_inst_min1_bfm (
		.sig_export (despertadorcpu_inst_min1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 despertadorcpu_inst_min2_bfm (
		.sig_export (despertadorcpu_inst_min2_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) despertadorcpu_inst_reset_bfm (
		.reset (despertadorcpu_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (despertadorcpu_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm despertadorcpu_inst_swinicio_bfm (
		.sig_export (despertadorcpu_inst_swinicio_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm despertadorcpu_inst_swmodo_bfm (
		.sig_export (despertadorcpu_inst_swmodo_bfm_conduit_export)  // conduit.export
	);

endmodule
