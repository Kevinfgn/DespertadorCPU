// DespertadorCPU.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DespertadorCPU (
		input  wire       btnapagar_export, // btnapagar.export
		input  wire       btnhora_export,   //   btnhora.export
		input  wire       btnmin_export,    //    btnmin.export
		output wire       buzzer_export,    //    buzzer.export
		input  wire       clk_clk,          //       clk.clk
		output wire [6:0] hora1_export,     //     hora1.export
		output wire [6:0] hora2_export,     //     hora2.export
		output wire [6:0] min1_export,      //      min1.export
		output wire [6:0] min2_export,      //      min2.export
		input  wire       reset_reset_n,    //     reset.reset_n
		input  wire       swinicio_export,  //  swinicio.export
		input  wire       swmodo_export     //    swmodo.export
	);

	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [13:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [13:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                      // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                        // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [9:0] mm_interconnect_0_memory_s1_address;                         // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                      // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                           // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                       // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                           // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_hora1_s1_chipselect;                       // mm_interconnect_0:hora1_s1_chipselect -> hora1:chipselect
	wire  [31:0] mm_interconnect_0_hora1_s1_readdata;                         // hora1:readdata -> mm_interconnect_0:hora1_s1_readdata
	wire   [1:0] mm_interconnect_0_hora1_s1_address;                          // mm_interconnect_0:hora1_s1_address -> hora1:address
	wire         mm_interconnect_0_hora1_s1_write;                            // mm_interconnect_0:hora1_s1_write -> hora1:write_n
	wire  [31:0] mm_interconnect_0_hora1_s1_writedata;                        // mm_interconnect_0:hora1_s1_writedata -> hora1:writedata
	wire         mm_interconnect_0_hora2_s1_chipselect;                       // mm_interconnect_0:hora2_s1_chipselect -> hora2:chipselect
	wire  [31:0] mm_interconnect_0_hora2_s1_readdata;                         // hora2:readdata -> mm_interconnect_0:hora2_s1_readdata
	wire   [1:0] mm_interconnect_0_hora2_s1_address;                          // mm_interconnect_0:hora2_s1_address -> hora2:address
	wire         mm_interconnect_0_hora2_s1_write;                            // mm_interconnect_0:hora2_s1_write -> hora2:write_n
	wire  [31:0] mm_interconnect_0_hora2_s1_writedata;                        // mm_interconnect_0:hora2_s1_writedata -> hora2:writedata
	wire         mm_interconnect_0_min1_s1_chipselect;                        // mm_interconnect_0:min1_s1_chipselect -> min1:chipselect
	wire  [31:0] mm_interconnect_0_min1_s1_readdata;                          // min1:readdata -> mm_interconnect_0:min1_s1_readdata
	wire   [1:0] mm_interconnect_0_min1_s1_address;                           // mm_interconnect_0:min1_s1_address -> min1:address
	wire         mm_interconnect_0_min1_s1_write;                             // mm_interconnect_0:min1_s1_write -> min1:write_n
	wire  [31:0] mm_interconnect_0_min1_s1_writedata;                         // mm_interconnect_0:min1_s1_writedata -> min1:writedata
	wire         mm_interconnect_0_min2_s1_chipselect;                        // mm_interconnect_0:min2_s1_chipselect -> min2:chipselect
	wire  [31:0] mm_interconnect_0_min2_s1_readdata;                          // min2:readdata -> mm_interconnect_0:min2_s1_readdata
	wire   [1:0] mm_interconnect_0_min2_s1_address;                           // mm_interconnect_0:min2_s1_address -> min2:address
	wire         mm_interconnect_0_min2_s1_write;                             // mm_interconnect_0:min2_s1_write -> min2:write_n
	wire  [31:0] mm_interconnect_0_min2_s1_writedata;                         // mm_interconnect_0:min2_s1_writedata -> min2:writedata
	wire  [31:0] mm_interconnect_0_btnhora_s1_readdata;                       // btnhora:readdata -> mm_interconnect_0:btnhora_s1_readdata
	wire   [1:0] mm_interconnect_0_btnhora_s1_address;                        // mm_interconnect_0:btnhora_s1_address -> btnhora:address
	wire  [31:0] mm_interconnect_0_btnmin_s1_readdata;                        // btnmin:readdata -> mm_interconnect_0:btnmin_s1_readdata
	wire   [1:0] mm_interconnect_0_btnmin_s1_address;                         // mm_interconnect_0:btnmin_s1_address -> btnmin:address
	wire  [31:0] mm_interconnect_0_btnapagar_s1_readdata;                     // btnapagar:readdata -> mm_interconnect_0:btnapagar_s1_readdata
	wire   [1:0] mm_interconnect_0_btnapagar_s1_address;                      // mm_interconnect_0:btnapagar_s1_address -> btnapagar:address
	wire  [31:0] mm_interconnect_0_swmodo_s1_readdata;                        // swmodo:readdata -> mm_interconnect_0:swmodo_s1_readdata
	wire   [1:0] mm_interconnect_0_swmodo_s1_address;                         // mm_interconnect_0:swmodo_s1_address -> swmodo:address
	wire         mm_interconnect_0_buzzer_s1_chipselect;                      // mm_interconnect_0:buzzer_s1_chipselect -> buzzer:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                        // buzzer:readdata -> mm_interconnect_0:buzzer_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                         // mm_interconnect_0:buzzer_s1_address -> buzzer:address
	wire         mm_interconnect_0_buzzer_s1_write;                           // mm_interconnect_0:buzzer_s1_write -> buzzer:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                       // mm_interconnect_0:buzzer_s1_writedata -> buzzer:writedata
	wire  [31:0] mm_interconnect_0_swinicio_s1_readdata;                      // swinicio:readdata -> mm_interconnect_0:swinicio_s1_readdata
	wire   [1:0] mm_interconnect_0_swinicio_s1_address;                       // mm_interconnect_0:swinicio_s1_address -> swinicio:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [btnapagar:reset_n, btnhora:reset_n, btnmin:reset_n, buzzer:reset_n, cpu:reset_n, hora1:reset_n, hora2:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, memory:reset, min1:reset_n, min2:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, swinicio:reset_n, swmodo:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, memory:reset_req, rst_translator:reset_req_in]

	DespertadorCPU_btnapagar btnapagar (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_btnapagar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_btnapagar_s1_readdata), //                    .readdata
		.in_port  (btnapagar_export)                         // external_connection.export
	);

	DespertadorCPU_btnapagar btnhora (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_btnhora_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_btnhora_s1_readdata), //                    .readdata
		.in_port  (btnhora_export)                         // external_connection.export
	);

	DespertadorCPU_btnapagar btnmin (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_btnmin_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_btnmin_s1_readdata), //                    .readdata
		.in_port  (btnmin_export)                         // external_connection.export
	);

	DespertadorCPU_buzzer buzzer (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                           // external_connection.export
	);

	DespertadorCPU_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DespertadorCPU_hora1 hora1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hora1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hora1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hora1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hora1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hora1_s1_readdata),   //                    .readdata
		.out_port   (hora1_export)                           // external_connection.export
	);

	DespertadorCPU_hora1 hora2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hora2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hora2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hora2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hora2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hora2_s1_readdata),   //                    .readdata
		.out_port   (hora2_export)                           // external_connection.export
	);

	DespertadorCPU_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	DespertadorCPU_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	DespertadorCPU_hora1 min1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_min1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_min1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_min1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_min1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_min1_s1_readdata),   //                    .readdata
		.out_port   (min1_export)                           // external_connection.export
	);

	DespertadorCPU_hora1 min2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_min2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_min2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_min2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_min2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_min2_s1_readdata),   //                    .readdata
		.out_port   (min2_export)                           // external_connection.export
	);

	DespertadorCPU_btnapagar swinicio (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_swinicio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_swinicio_s1_readdata), //                    .readdata
		.in_port  (swinicio_export)                         // external_connection.export
	);

	DespertadorCPU_btnapagar swmodo (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_swmodo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_swmodo_s1_readdata), //                    .readdata
		.in_port  (swmodo_export)                         // external_connection.export
	);

	DespertadorCPU_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	DespertadorCPU_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                              // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                   (cpu_data_master_address),                                     //                 cpu_data_master.address
		.cpu_data_master_waitrequest               (cpu_data_master_waitrequest),                                 //                                .waitrequest
		.cpu_data_master_byteenable                (cpu_data_master_byteenable),                                  //                                .byteenable
		.cpu_data_master_read                      (cpu_data_master_read),                                        //                                .read
		.cpu_data_master_readdata                  (cpu_data_master_readdata),                                    //                                .readdata
		.cpu_data_master_write                     (cpu_data_master_write),                                       //                                .write
		.cpu_data_master_writedata                 (cpu_data_master_writedata),                                   //                                .writedata
		.cpu_data_master_debugaccess               (cpu_data_master_debugaccess),                                 //                                .debugaccess
		.cpu_instruction_master_address            (cpu_instruction_master_address),                              //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest        (cpu_instruction_master_waitrequest),                          //                                .waitrequest
		.cpu_instruction_master_read               (cpu_instruction_master_read),                                 //                                .read
		.cpu_instruction_master_readdata           (cpu_instruction_master_readdata),                             //                                .readdata
		.btnapagar_s1_address                      (mm_interconnect_0_btnapagar_s1_address),                      //                    btnapagar_s1.address
		.btnapagar_s1_readdata                     (mm_interconnect_0_btnapagar_s1_readdata),                     //                                .readdata
		.btnhora_s1_address                        (mm_interconnect_0_btnhora_s1_address),                        //                      btnhora_s1.address
		.btnhora_s1_readdata                       (mm_interconnect_0_btnhora_s1_readdata),                       //                                .readdata
		.btnmin_s1_address                         (mm_interconnect_0_btnmin_s1_address),                         //                       btnmin_s1.address
		.btnmin_s1_readdata                        (mm_interconnect_0_btnmin_s1_readdata),                        //                                .readdata
		.buzzer_s1_address                         (mm_interconnect_0_buzzer_s1_address),                         //                       buzzer_s1.address
		.buzzer_s1_write                           (mm_interconnect_0_buzzer_s1_write),                           //                                .write
		.buzzer_s1_readdata                        (mm_interconnect_0_buzzer_s1_readdata),                        //                                .readdata
		.buzzer_s1_writedata                       (mm_interconnect_0_buzzer_s1_writedata),                       //                                .writedata
		.buzzer_s1_chipselect                      (mm_interconnect_0_buzzer_s1_chipselect),                      //                                .chipselect
		.cpu_debug_mem_slave_address               (mm_interconnect_0_cpu_debug_mem_slave_address),               //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                 (mm_interconnect_0_cpu_debug_mem_slave_write),                 //                                .write
		.cpu_debug_mem_slave_read                  (mm_interconnect_0_cpu_debug_mem_slave_read),                  //                                .read
		.cpu_debug_mem_slave_readdata              (mm_interconnect_0_cpu_debug_mem_slave_readdata),              //                                .readdata
		.cpu_debug_mem_slave_writedata             (mm_interconnect_0_cpu_debug_mem_slave_writedata),             //                                .writedata
		.cpu_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_debug_mem_slave_byteenable),            //                                .byteenable
		.cpu_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),           //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),           //                                .debugaccess
		.hora1_s1_address                          (mm_interconnect_0_hora1_s1_address),                          //                        hora1_s1.address
		.hora1_s1_write                            (mm_interconnect_0_hora1_s1_write),                            //                                .write
		.hora1_s1_readdata                         (mm_interconnect_0_hora1_s1_readdata),                         //                                .readdata
		.hora1_s1_writedata                        (mm_interconnect_0_hora1_s1_writedata),                        //                                .writedata
		.hora1_s1_chipselect                       (mm_interconnect_0_hora1_s1_chipselect),                       //                                .chipselect
		.hora2_s1_address                          (mm_interconnect_0_hora2_s1_address),                          //                        hora2_s1.address
		.hora2_s1_write                            (mm_interconnect_0_hora2_s1_write),                            //                                .write
		.hora2_s1_readdata                         (mm_interconnect_0_hora2_s1_readdata),                         //                                .readdata
		.hora2_s1_writedata                        (mm_interconnect_0_hora2_s1_writedata),                        //                                .writedata
		.hora2_s1_chipselect                       (mm_interconnect_0_hora2_s1_chipselect),                       //                                .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                .chipselect
		.memory_s1_address                         (mm_interconnect_0_memory_s1_address),                         //                       memory_s1.address
		.memory_s1_write                           (mm_interconnect_0_memory_s1_write),                           //                                .write
		.memory_s1_readdata                        (mm_interconnect_0_memory_s1_readdata),                        //                                .readdata
		.memory_s1_writedata                       (mm_interconnect_0_memory_s1_writedata),                       //                                .writedata
		.memory_s1_byteenable                      (mm_interconnect_0_memory_s1_byteenable),                      //                                .byteenable
		.memory_s1_chipselect                      (mm_interconnect_0_memory_s1_chipselect),                      //                                .chipselect
		.memory_s1_clken                           (mm_interconnect_0_memory_s1_clken),                           //                                .clken
		.min1_s1_address                           (mm_interconnect_0_min1_s1_address),                           //                         min1_s1.address
		.min1_s1_write                             (mm_interconnect_0_min1_s1_write),                             //                                .write
		.min1_s1_readdata                          (mm_interconnect_0_min1_s1_readdata),                          //                                .readdata
		.min1_s1_writedata                         (mm_interconnect_0_min1_s1_writedata),                         //                                .writedata
		.min1_s1_chipselect                        (mm_interconnect_0_min1_s1_chipselect),                        //                                .chipselect
		.min2_s1_address                           (mm_interconnect_0_min2_s1_address),                           //                         min2_s1.address
		.min2_s1_write                             (mm_interconnect_0_min2_s1_write),                             //                                .write
		.min2_s1_readdata                          (mm_interconnect_0_min2_s1_readdata),                          //                                .readdata
		.min2_s1_writedata                         (mm_interconnect_0_min2_s1_writedata),                         //                                .writedata
		.min2_s1_chipselect                        (mm_interconnect_0_min2_s1_chipselect),                        //                                .chipselect
		.swinicio_s1_address                       (mm_interconnect_0_swinicio_s1_address),                       //                     swinicio_s1.address
		.swinicio_s1_readdata                      (mm_interconnect_0_swinicio_s1_readdata),                      //                                .readdata
		.swmodo_s1_address                         (mm_interconnect_0_swmodo_s1_address),                         //                       swmodo_s1.address
		.swmodo_s1_readdata                        (mm_interconnect_0_swmodo_s1_readdata),                        //                                .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                      timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                .chipselect
	);

	DespertadorCPU_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
